module top_neurex (
  input clk,
  input rstn,
  input 
